module arrays();

    wire [7 : 0] vect;
    
    wire arr[3 : 0];
    
    wire [7 : 0] arr_vec[3 : 0];
    
    
endmodule